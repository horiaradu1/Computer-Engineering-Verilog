//Verilog HDL for "MU0_lib", "mux_2to1_12bit" "functional"


module mux_2to1_12bit ( output reg [11:0] q,
			input [11:0] a,
			input [11:0] b,
			input sel );

endmodule
