// Verilog stimulus file.
// Please do not create a module in this file.
/*

#VALUE      creates a delay of VALUE ns
a=VALUE;    sets the value of input 'a' to VALUE
$stop;      tells the simulator to stop

*/

initial
begin
#100 bcd=0;

// Enter you stimulus below this line
// Make sure you test all input combinations with a delay
// -------------------------------------------------------





// -------------------------------------------------------
// Please make sure your stimulus is above this line
 
#100 $stop;
end
