// Verilog HDL for "COMP12111_lib", "sevensegmentdecoder" "functional"
// Created P W Nutter, 20/3/19
//
// Add your comments here ...


module sevensegmentdecoder (input [3:0] bcd,
			    output reg 	[7:0] segments);

// create an always block to represent the desired behaviour of the
// combinatorial design
// -----------------------------------------------------------------







endmodule  // end of module sevensegmentdecoder
