//Verilog HDL for "TEST", "fulladder" "functional"


module fulladder ( );

endmodule
